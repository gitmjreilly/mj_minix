library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
library UNISIM;
use UNISIM.VComponents.all;

entity video_card is
   Port ( addr_bus : in  STD_LOGIC_VECTOR (11 downto 0);
           data_bus : inout  STD_LOGIC_VECTOR (15 downto 0);
           n_wr : in  STD_LOGIC;
           n_rd : in  STD_LOGIC;
           n_cs : in  STD_LOGIC;
           clock : in  STD_LOGIC;

	 			reset : in std_logic;
				r_out : out std_logic;
				g_out : out std_logic;
				b_out : out std_logic;
				hsyncb : out std_logic;
           	vsyncb : out std_logic);
end video_card;

architecture Behavioral of video_card is

	constant max_h_count : integer := 793;
	constant min_h_pulse_count : integer := 653;
	constant max_h_pulse_count : integer := 748;

	constant max_v_count : integer := 527;
	constant min_v_pulse_count : integer := 490;
	constant max_v_pulse_count : integer := 492;

--	constant max_v_count : integer := 627;
--	constant min_v_pulse_count : integer := 590;
--	constant max_v_pulse_count : integer := 592;


	signal h_sync_internal : std_logic;
	signal h_count : std_logic_vector(9 downto 0);
	signal v_count : std_logic_vector(8 downto 0);
	signal clock_counter : std_logic_vector(1 downto 0);
	signal video_clock : std_logic;
	signal VERTICAL_OFFSET_ADDR : std_logic_vector(7 downto 0);
	signal HORIZONTAL_OFFSET_ADDR : std_logic_vector(7 downto 0);
	signal video_out : std_logic;

	signal data_word_16 : std_logic_vector(15 downto 0);
	signal word_number : std_logic_vector(5 downto 0);
	signal video_buffer : std_logic_vector(639 downto 0);
	signal VIDEO_DATA_OUT : STD_LOGIC_VECTOR(0 downto 0);      -- 1-bit Data Output
	signal VIDEO_DATA_OUT_0 : STD_LOGIC_VECTOR(0 downto 0);
	signal VIDEO_DATA_OUT_1 : STD_LOGIC_VECTOR(0 downto 0);
	signal VIDEO_DATA_OUT_2 : STD_LOGIC_VECTOR(0 downto 0);
	signal VIDEO_DATA_OUT_3 : STD_LOGIC_VECTOR(0 downto 0);
   signal CONSTRUCTED_VIDEO_ADDR : STD_LOGIC_VECTOR(15 downto 0);

	signal CPU_DATA_OUT : STD_LOGIC_VECTOR(15 downto 0);
	signal CPU_DATA_OUT_0 : STD_LOGIC_VECTOR(15 downto 0);
	signal CPU_DATA_OUT_1 : STD_LOGIC_VECTOR(15 downto 0);
	signal CPU_DATA_OUT_2 : STD_LOGIC_VECTOR(15 downto 0);
	signal CPU_DATA_OUT_3 : STD_LOGIC_VECTOR(15 downto 0);
	signal PADDED_ADDR : STD_LOGIC_VECTOR(9 downto 0);
	signal OUTPUT_ENABLE : STD_LOGIC;
	signal DOPB : STD_LOGIC_VECTOR(1 downto 0);

	signal UPPER_2_VIDEO_ADDRESS_BITS : STD_LOGIC_VECTOR(1 DOWNTO 0);
	signal UPPER_2_CPU_ADDRESS_BITS : STD_LOGIC_VECTOR(1 DOWNTO 0);
	
	signal RAM_CPU_ENABLE_0 : STD_LOGIC;
	signal RAM_CPU_ENABLE_1 : STD_LOGIC;
	signal RAM_CPU_ENABLE_2 : STD_LOGIC;
	signal RAM_CPU_ENABLE_3 : STD_LOGIC;


begin

  RAMB16_S1_S18_inst_0 : RAMB16_S1_S18
   generic map (
      INIT_A => X"0", --  Value of output RAM registers on Port A at startup
      INIT_B => X"00000", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"0", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"00000", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "READ_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL" 
      -- The following INIT_xx declarations specify the initial contents of the RAM
      -- Port A Address 0 to 4095, Port B Address 0 to 255
      INIT_00 => X"FFFFFFFFFFFFFFFFFFFFF00000000000000000000000FFFFFFFFFFFFFFFFFFF0",
      INIT_01 => X"0000011111111111111110000000000000000000000011111111111111111111",
      INIT_02 => X"3333333333333333333300000000000000000000000033333333333333333333",
      INIT_03 => X"7777777777777777770000000000000000000000000777777777777777777777",
      INIT_04 => X"FFFFFFFFFFFFFFFFFFFFF0000000000000000000000FFFFFFFFFFFFFFFFFFFFF",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 4096 to 8191, Port B Address 256 to 511
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000FFF000000000000000000000000000000000000",
      INIT_12 => X"000000000000000000000F0FF0000F0F00000000000000000000000000000000",
      INIT_13 => X"0000000000000000000FF00000000000F0000000000000000000000000000000",
      INIT_14 => X"000000000000000000F00000000000000F000000000000000000000000000000",
      INIT_15 => X"00000000000000000F0000000000000000F00000000000000000000000000000",
      INIT_16 => X"00000000000000F0F000000000000000000F0000000000000000000000000000",
      INIT_17 => X"0000000000000F0000000000000000000000F000000000000000000000000000",
      INIT_18 => X"0000000000000FF0000000000000000000000F00000000000000000000000000",
      INIT_19 => X"000000000000000F0000000000000000000000F0000000000000000000000000",
      INIT_1A => X"0000000000000000F00000000000000000000F0F000000000000000000000000",
      INIT_1B => X"00000000000000000FFF00000000000FFF0F0000000000000000000000000000",
      INIT_1C => X"0000000000000000000F00000000FFF000000000000000000000000000000000",
      INIT_1D => X"000000000000000000F0F000000F000000000000000000000000000000000000",
      INIT_1E => X"000000000000000000000F0000F0000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000FFFF00000000000000000000000000000000000000",
      -- Port A Address 8192 to 12287, Port B Address 512 to 767
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 12288 to 16383, Port B Address 768 to 1023
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- The next set of INITP_xx are for the parity bits
      -- Port B Address 0 to 255
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port B Address 256 to 511
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port B Address 512 to 767
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port B Address 768 to 1023 
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => VIDEO_DATA_OUT_0,      -- Port A 1-bit Data Output
      DOB => CPU_DATA_OUT_0,       -- Port B 16-bit Data Output
--      DOPB => DOPB,     -- Port B 2-bit Parity Output
      ADDRA => CONSTRUCTED_VIDEO_ADDR(13 downto 0),   -- 14-bit Address (created by video circuit)
      ADDRB => PADDED_ADDR,   -- Port B 10-bit Address Input
      CLKA => (NOT CLOCK),     -- Port A Clock
      CLKB => (NOT CLOCK),     -- Port B Clock
      DIA => "1",       -- Port A Input - NOT used Port A is READ ONLY by Vid circuit
      DIB => DATA_BUS,       -- Port B 16-bit Data Input
      DIPB => "00",     -- Port-B 2-bit parity Input
      ENA => '1',       -- Port A RAM Enable Input
      ENB => RAM_CPU_ENABLE_0,     -- PortB RAM Enable Input
      SSRA => '0',     -- Port A Synchronous Set/Reset Input
      SSRB => '0',     -- Port B Synchronous Set/Reset Input
      WEA => '0',       -- Port A Write Enable Input
      WEB => (NOT N_WR)        -- Port B Write Enable Input
   );

  RAMB16_S1_S18_inst_1 : RAMB16_S1_S18
   generic map (
      INIT_A => X"0", --  Value of output RAM registers on Port A at startup
      INIT_B => X"00000", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"0", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"00000", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "READ_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL" 
      -- The following INIT_xx declarations specify the initial contents of the RAM
      -- Port A Address 0 to 4095, Port B Address 0 to 255
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 4096 to 8191, Port B Address 256 to 511
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000F00000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000F00000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000F00000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000F00000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000F00000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000F00000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000F00000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000F00000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000F00000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000F00000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000F00000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000F00000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000F00000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000F00000000000000000000000000000000000000",
      -- Port A Address 8192 to 12287, Port B Address 512 to 767
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 12288 to 16383, Port B Address 768 to 1023
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- The next set of INITP_xx are for the parity bits
      -- Port B Address 0 to 255
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port B Address 256 to 511
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port B Address 512 to 767
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port B Address 768 to 1023 
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => VIDEO_DATA_OUT_1,      -- Port A 1-bit Data Output
      DOB => CPU_DATA_OUT_1,       -- Port B 16-bit Data Output
--      DOPB => DOPB,     -- Port B 2-bit Parity Output
      ADDRA => CONSTRUCTED_VIDEO_ADDR(13 downto 0),   -- 14-bit Address (created by video circuit)
      ADDRB => PADDED_ADDR,   -- Port B 10-bit Address Input
      CLKA => (NOT CLOCK),     -- Port A Clock
      CLKB => (NOT CLOCK),     -- Port B Clock
      DIA => "1",       -- Port A Input - NOT used Port A is READ ONLY by Vid circuit
      DIB => DATA_BUS,       -- Port B 16-bit Data Input
      DIPB => "00",     -- Port-B 2-bit parity Input
      ENA => '1',       -- Port A RAM Enable Input
      ENB => RAM_CPU_ENABLE_1,     -- PortB RAM Enable Input
      SSRA => '0',     -- Port A Synchronous Set/Reset Input
      SSRB => '0',     -- Port B Synchronous Set/Reset Input
      WEA => '0',       -- Port A Write Enable Input
      WEB => (NOT N_WR)        -- Port B Write Enable Input
   );

  RAMB16_S1_S18_inst_2 : RAMB16_S1_S18
   generic map (
      INIT_A => X"0", --  Value of output RAM registers on Port A at startup
      INIT_B => X"00000", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"0", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"00000", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "READ_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL" 
      -- The following INIT_xx declarations specify the initial contents of the RAM
      -- Port A Address 0 to 4095, Port B Address 0 to 255
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 4096 to 8191, Port B Address 256 to 511
      INIT_10 => X"0000000000000000000F000000000000000000000F0000000000000000000000",
      INIT_11 => X"0000000000000000000F000000000000000000000F0000000000000000000000",
      INIT_12 => X"0000000000000000000F000000000000000000000F0000000000000000000000",
      INIT_13 => X"0000000000000000000F000000000000000000000F0000000000000000000000",
      INIT_14 => X"0000000000000000000F000000000000000000000F0000000000000000000000",
      INIT_15 => X"0000000000000000000F000000000000000000000F0000000000000000000000",
      INIT_16 => X"0000000000000000000F000000000000000000000F0000000000000000000000",
      INIT_17 => X"0000000000000000000F000000000000000000000F0000000000000000000000",
      INIT_18 => X"0000000000000000000F000000000000000000000F0000000000000000000000",
      INIT_19 => X"0000000000000000000F000000000000000000000F0000000000000000000000",
      INIT_1A => X"0000000000000000000F000000000000000000000F0000000000000000000000",
      INIT_1B => X"0000000000000000000F000000000000000000000F0000000000000000000000",
      INIT_1C => X"0000000000000000000F000000000000000000000F0000000000000000000000",
      INIT_1D => X"0000000000000000000F000000000000000000000F0000000000000000000000",
      INIT_1E => X"0000000000000000000F000000000000000000000F0000000000000000000000",
      INIT_1F => X"0000000000000000000F00000000000000000000000000000000000000000000",
      -- Port A Address 8192 to 12287, Port B Address 512 to 767
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 12288 to 16383, Port B Address 768 to 1023
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- The next set of INITP_xx are for the parity bits
      -- Port B Address 0 to 255
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port B Address 256 to 511
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port B Address 512 to 767
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port B Address 768 to 1023 
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => VIDEO_DATA_OUT_2,      -- Port A 1-bit Data Output
      DOB => CPU_DATA_OUT_2,       -- Port B 16-bit Data Output
--      DOPB => DOPB,     -- Port B 2-bit Parity Output
      ADDRA => CONSTRUCTED_VIDEO_ADDR(13 downto 0),   -- 14-bit Address (created by video circuit)
      ADDRB => PADDED_ADDR,   -- Port B 10-bit Address Input
      CLKA => (NOT CLOCK),     -- Port A Clock
      CLKB => (NOT CLOCK),     -- Port B Clock
      DIA => "1",       -- Port A Input - NOT used Port A is READ ONLY by Vid circuit
      DIB => DATA_BUS,       -- Port B 16-bit Data Input
      DIPB => "00",     -- Port-B 2-bit parity Input
      ENA => '1',       -- Port A RAM Enable Input
      ENB => RAM_CPU_ENABLE_2,     -- PortB RAM Enable Input
      SSRA => '0',     -- Port A Synchronous Set/Reset Input
      SSRB => '0',     -- Port B Synchronous Set/Reset Input
      WEA => '0',       -- Port A Write Enable Input
      WEB => (NOT N_WR)        -- Port B Write Enable Input
   );

  RAMB16_S1_S18_inst_3 : RAMB16_S1_S18
   generic map (
      INIT_A => X"0", --  Value of output RAM registers on Port A at startup
      INIT_B => X"00000", --  Value of output RAM registers on Port B at startup
      SRVAL_A => X"0", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"00000", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "WRITE_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "READ_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL" 
      -- The following INIT_xx declarations specify the initial contents of the RAM
      -- Port A Address 0 to 4095, Port B Address 0 to 255
      INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 4096 to 8191, Port B Address 256 to 511
      INIT_10 => X"000000000000000F00000000000000000000F000000000000000F00000000000",
      INIT_11 => X"000000000000000F00000000000000000000F000000000000000F00000000000",
      INIT_12 => X"000000000000000F00000000000000000000FF00000000000000F00000000000",
      INIT_13 => X"000000000000000F00000000000000000000F000000000000000F00000000000",
      INIT_14 => X"000000000000000F00000000000000000000F000000000000000F00000000000",
      INIT_15 => X"000000000000000F00000000000000000000F000000000000000F00000000000",
      INIT_16 => X"000000000000000F00000000000000000000F000000000000000F00000000000",
      INIT_17 => X"000000000000000F00000000000000000000F000000000000000F00000000000",
      INIT_18 => X"000000000000000F00000000000000000000F000000000000000F00000000000",
      INIT_19 => X"000000000000000F00000000000000000000F000000000000000F00000000000",
      INIT_1A => X"000000000000000F00000000000000000000F000000000000000F00000000000",
      INIT_1B => X"000000000000000F00000000000000000000F000000000000000F00000000000",
      INIT_1C => X"000000000000000F00000000000000000000F000000000000000F00000000000",
      INIT_1D => X"000000000000000F00000000000000000000F000000000000000F00000000000",
      INIT_1E => X"000000000000000F00000000000000000000F000000000000000F00000000000",
      INIT_1F => X"000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000",
      -- Port A Address 8192 to 12287, Port B Address 512 to 767
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 12288 to 16383, Port B Address 768 to 1023
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"00000000000000000000F0F0F0F0F0F0F0F0F0F0F00000000000000000000000",
      INIT_3F => X"00000000000000000000AAAAAAAAAAAAAAAAAAAAA00000000000000000000000",
      -- The next set of INITP_xx are for the parity bits
      -- Port B Address 0 to 255
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port B Address 256 to 511
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port B Address 512 to 767
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port B Address 768 to 1023 
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => VIDEO_DATA_OUT_3,     -- Port A 1-bit Data Output
      DOB => CPU_DATA_OUT_3,       -- Port B 16-bit Data Output
--      DOPB => DOPB,     -- Port B 2-bit Parity Output
      ADDRA => CONSTRUCTED_VIDEO_ADDR(13 downto 0),   -- 14-bit Address (created by video circuit)
      ADDRB => PADDED_ADDR,   -- Port B 10-bit Address Input
      CLKA => (NOT CLOCK),     -- Port A Clock
      CLKB => (NOT CLOCK),     -- Port B Clock
      DIA => "1",       -- Port A Input - NOT used Port A is READ ONLY by Vid circuit
      DIB => DATA_BUS,       -- Port B 16-bit Data Input
      DIPB => "00",     -- Port-B 2-bit parity Input
      ENA => '1',       -- Port A RAM Enable Input
      ENB => RAM_CPU_ENABLE_3,     -- PortB RAM Enable Input
      SSRA => '0',     -- Port A Synchronous Set/Reset Input
      SSRB => '0',     -- Port B Synchronous Set/Reset Input
      WEA => '0',       -- Port A Write Enable Input
      WEB => (NOT N_WR)        -- Port B Write Enable Input
   );

	UPPER_2_CPU_ADDRESS_BITS <= ADDR_BUS(11 DOWNTO 10);
	PADDED_ADDR <= ADDR_BUS(9 DOWNTO 0);

	output_enable <= (n_wr) and (NOT n_cs);
	

	CPU_DATA_OUT <= 
		CPU_DATA_OUT_0 WHEN UPPER_2_CPU_ADDRESS_BITS = "00" ELSE
		CPU_DATA_OUT_1 WHEN UPPER_2_CPU_ADDRESS_BITS = "01" ELSE
		CPU_DATA_OUT_2 WHEN UPPER_2_CPU_ADDRESS_BITS = "10" ELSE
		CPU_DATA_OUT_3 WHEN UPPER_2_CPU_ADDRESS_BITS = "11";

	data_bus <= CPU_DATA_OUT when (output_enable = '1') else "ZZZZZZZZZZZZZZZZ";



	hsyncb <= h_sync_internal;

	clock_counter_proc : process(clock, reset) 
	begin
		if (reset = '1') then
			clock_counter <= (others => '0');
		elsif (rising_edge(clock)) then
			clock_counter <= clock_counter + 1;
		end if;
	end process;

--	video_clock <= clock_counter(0);
	video_clock <= clock;

	--
	-- Horizontal Pixel Counter
	--
	h_pixel_clock: process (video_clock, reset)
	begin
		if (reset = '1') then
			h_count <= (others => '0');
		elsif (rising_edge(video_clock)) then
			if (h_count < max_h_count) then
				h_count <= h_count + 1;
			else
				h_count <= (others => '0');
			end if;
		end if;
	end process;

	--
	-- Horizontal Sync Pulse
	--
	h_sync_proc: process (video_clock, reset)
	begin
		if (reset = '1') then
			h_sync_internal <= '1';
		elsif (rising_edge(video_clock)) then
			if (h_count >= min_h_pulse_count and h_count < max_h_pulse_count) then
				h_sync_internal <= '0';
			else
				h_sync_internal <= '1';
			end if;
		end if;
	end process	;

	--
	-- Vertical Line Counter (uses horizontal sync pulse)
	v_line_counter: process (h_sync_internal, reset)
	begin
		if (reset = '1') then
			v_count <= (others => '0');
		elsif (rising_edge(h_sync_internal)) then
			if (v_count < max_v_count) then
				v_count <= v_count + 1;
			else
				v_count <= (others => '0');
			end if;
		end if;
	end process;

	--
	-- Vertical Sync Pulse Generator
	--
	v_sync_proc: process (h_sync_internal, reset)
	begin
		if (reset = '1') then
			vsyncb <= '1';
		elsif (rising_edge(h_sync_internal)) then
			if (v_count >= min_v_pulse_count and v_count < max_v_pulse_count) then
				vsyncb <= '0';
			else
				vsyncb <= '1';
			end if;
		end if;
	end process;


	VERTICAL_OFFSET_ADDR <= v_count(7 downto 0) - "01110000"; -- (480 - 256)/2 = 112
	HORIZONTAL_OFFSET_ADDR <= h_count(7 downto 0) - "11000000"; -- (640-256)/2 = 192
	CONSTRUCTED_VIDEO_ADDR <= VERTICAL_OFFSET_ADDR & HORIZONTAL_OFFSET_ADDR(7 downto 0);
	UPPER_2_VIDEO_ADDRESS_BITS <= CONSTRUCTED_VIDEO_ADDR(15 DOWNTO 14);

	VIDEO_DATA_OUT <= 
		VIDEO_DATA_OUT_0 WHEN UPPER_2_VIDEO_ADDRESS_BITS = "00" ELSE
		VIDEO_DATA_OUT_1 WHEN UPPER_2_VIDEO_ADDRESS_BITS = "01" ELSE
		VIDEO_DATA_OUT_2 WHEN UPPER_2_VIDEO_ADDRESS_BITS = "10" ELSE
		VIDEO_DATA_OUT_3 WHEN UPPER_2_VIDEO_ADDRESS_BITS = "11";

	RAM_CPU_ENABLE_0 <= (NOT N_CS) WHEN UPPER_2_CPU_ADDRESS_BITS = "00" ELSE '0';
	RAM_CPU_ENABLE_1 <= (NOT N_CS) WHEN UPPER_2_CPU_ADDRESS_BITS = "01" ELSE '0';
	RAM_CPU_ENABLE_2 <= (NOT N_CS) WHEN UPPER_2_CPU_ADDRESS_BITS = "10" ELSE '0';
	RAM_CPU_ENABLE_3 <= (NOT N_CS) WHEN UPPER_2_CPU_ADDRESS_BITS = "11" ELSE '0';

	--
	-- Process to draw a box on the screen
	--
	draw_proc : process (video_clock)
	begin
		if (	(h_count >= 192 and h_count < (256 + 192))  and
				(v_count >= 112 and v_count < (256+112) ) ) then
				video_out <= VIDEO_DATA_OUT(0);
		else
				video_out <= '0';
		end if;
	end process;





	r_out <= '0';
	g_out <= video_out;
	b_out <= '0';
		

end Behavioral;
