library IEEE; 

use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity rom is
    Port ( addr : in std_logic_vector(15 downto 0);
           data : out std_logic_vector(15 downto 0);
           cs : in std_logic);
end rom;


architecture Behavioral of rom is

  signal output : std_logic_vector(15 downto 0);

begin
   output <= 
--
--x"0002" when (addr =  x"0") else
--x"0017" when (addr =  x"1") else
--x"0002" when (addr =  x"2") else
--x"0002" when (addr =  x"3") else
--x"0018" when (addr =  x"4") else
--x"0003" when (addr =  x"5") else
--

-- Pat's Original
x"000A" when (addr =  x"0") else
x"006F" when (addr =  x"1") else
x"0002" when (addr =  x"2") else
x"F001" when (addr =  x"3") else
x"0009" when (addr =  x"4") else
x"0002" when (addr =  x"5") else

x"0001" when (addr =  x"6") else
x"001B" when (addr =  x"7") else
x"0002" when (addr =  x"8") else
x"0001" when (addr =  x"9") else
x"001F" when (addr =  x"a") else
x"000C" when (addr =  x"b") else
x"0002" when (addr =  x"c") else
x"0002" when (addr =  x"d") else
x"F000" when (addr =  x"e") else
x"0008" when (addr =  x"f") else
x"000B" when (addr =  x"10") else
x"0002" when (addr =  x"11") else
x"F001" when (addr =  x"12") else
x"0009" when (addr =  x"13") else
x"0002" when (addr =  x"14") else
x"0002" when (addr =  x"15") else
x"001B" when (addr =  x"16") else
x"0002" when (addr =  x"17") else
x"0002" when (addr =  x"18") else
x"001F" when (addr =  x"19") else
x"000C" when (addr =  x"1a") else
x"0011" when (addr =  x"1b") else
x"000B" when (addr =  x"1c") else
x"000A" when (addr =  x"1d") else
x"0011" when (addr =  x"1e") else
x"0002" when (addr =  x"1f") else
x"F000" when (addr =  x"20") else
x"0009" when (addr =  x"21") else
x"000B" when (addr =  x"22") else
x"0015" when (addr =  x"23") else
x"0019" when (addr =  x"24") else
x"001A" when (addr =  x"25") else
x"000B" when (addr =  x"26") else
x"000A" when (addr =  x"27") else
x"001D" when (addr =  x"28") else
x"0013" when (addr =  x"29") else
x"0002" when (addr =  x"2a") else
x"0040" when (addr =  x"2b") else
x"0005" when (addr =  x"2c") else
x"000C" when (addr =  x"2d") else
x"0033" when (addr =  x"2e") else
x"0002" when (addr =  x"2f") else
x"0030" when (addr =  x"30") else
x"0004" when (addr =  x"31") else
x"0035" when (addr =  x"32") else
x"0002" when (addr =  x"33") else
x"0037" when (addr =  x"34") else
x"0019" when (addr =  x"35") else
x"000B" when (addr =  x"36") else
x"000A" when (addr =  x"37") else
x"0027" when (addr =  x"38") else
x"0002" when (addr =  x"39") else
x"1000" when (addr =  x"3a") else
x"001E" when (addr =  x"3b") else
x"000A" when (addr =  x"3c") else
x"0027" when (addr =  x"3d") else
x"0002" when (addr =  x"3e") else
x"0100" when (addr =  x"3f") else
x"001E" when (addr =  x"40") else
x"0018" when (addr =  x"41") else
x"000A" when (addr =  x"42") else
x"0027" when (addr =  x"43") else
x"0002" when (addr =  x"44") else
x"0010" when (addr =  x"45") else
x"001E" when (addr =  x"46") else
x"0018" when (addr =  x"47") else
x"000A" when (addr =  x"48") else
x"0027" when (addr =  x"49") else
x"0018" when (addr =  x"4a") else
x"000B" when (addr =  x"4b") else
x"0002" when (addr =  x"4c") else
x"000D" when (addr =  x"4d") else
x"000A" when (addr =  x"4e") else
x"0002" when (addr =  x"4f") else
x"0002" when (addr =  x"50") else
x"000A" when (addr =  x"51") else
x"000A" when (addr =  x"52") else
x"0002" when (addr =  x"53") else
x"000B" when (addr =  x"54") else
x"0002" when (addr =  x"55") else
x"0058" when (addr =  x"56") else
x"000B" when (addr =  x"57") else
x"FFFF" when (addr =  x"58") else
x"000E" when (addr =  x"59") else
x"000E" when (addr =  x"5a") else
x"0013" when (addr =  x"5b") else
x"0002" when (addr =  x"5c") else
x"0000" when (addr =  x"5d") else
x"000A" when (addr =  x"5e") else
x"0023" when (addr =  x"5f") else
x"000C" when (addr =  x"60") else
x"0069" when (addr =  x"61") else
x"0002" when (addr =  x"62") else
x"0001" when (addr =  x"63") else
x"0019" when (addr =  x"64") else
x"000D" when (addr =  x"65") else
x"0009" when (addr =  x"66") else
x"000D" when (addr =  x"67") else
x"000B" when (addr =  x"68") else
x"0007" when (addr =  x"69") else
x"0002" when (addr =  x"6a") else
x"0001" when (addr =  x"6b") else
x"0018" when (addr =  x"6c") else
x"000D" when (addr =  x"6d") else
x"000B" when (addr =  x"6e") else
x"000A" when (addr =  x"6f") else
x"004C" when (addr =  x"70") else
x"000A" when (addr =  x"71") else
x"004C" when (addr =  x"72") else
x"0002" when (addr =  x"73") else
x"002D" when (addr =  x"74") else
x"000A" when (addr =  x"75") else
x"0002" when (addr =  x"76") else
x"0002" when (addr =  x"77") else
x"002D" when (addr =  x"78") else
x"000A" when (addr =  x"79") else
x"0002" when (addr =  x"7a") else
x"0002" when (addr =  x"7b") else
x"002D" when (addr =  x"7c") else
x"000A" when (addr =  x"7d") else
x"0002" when (addr =  x"7e") else
x"0002" when (addr =  x"7f") else
x"002D" when (addr =  x"80") else
x"000A" when (addr =  x"81") else
x"0002" when (addr =  x"82") else
x"0002" when (addr =  x"83") else
x"002D" when (addr =  x"84") else
x"000A" when (addr =  x"85") else
x"0002" when (addr =  x"86") else
x"0002" when (addr =  x"87") else
x"002D" when (addr =  x"88") else
x"000A" when (addr =  x"89") else
x"0002" when (addr =  x"8a") else
x"0002" when (addr =  x"8b") else
x"002D" when (addr =  x"8c") else
x"000A" when (addr =  x"8d") else
x"0002" when (addr =  x"8e") else
x"0002" when (addr =  x"8f") else
x"002D" when (addr =  x"90") else
x"000A" when (addr =  x"91") else
x"0002" when (addr =  x"92") else
x"0002" when (addr =  x"93") else
x"002D" when (addr =  x"94") else
x"000A" when (addr =  x"95") else
x"0002" when (addr =  x"96") else
x"0002" when (addr =  x"97") else
x"002D" when (addr =  x"98") else
x"000A" when (addr =  x"99") else
x"0002" when (addr =  x"9a") else
x"0002" when (addr =  x"9b") else
x"002D" when (addr =  x"9c") else
x"000A" when (addr =  x"9d") else
x"0002" when (addr =  x"9e") else
x"0002" when (addr =  x"9f") else
x"002D" when (addr =  x"a0") else
x"000A" when (addr =  x"a1") else
x"0002" when (addr =  x"a2") else
x"0002" when (addr =  x"a3") else
x"002D" when (addr =  x"a4") else
x"000A" when (addr =  x"a5") else
x"0002" when (addr =  x"a6") else
x"0002" when (addr =  x"a7") else
x"002D" when (addr =  x"a8") else
x"000A" when (addr =  x"a9") else
x"0002" when (addr =  x"aa") else
x"0002" when (addr =  x"ab") else
x"002D" when (addr =  x"ac") else
x"000A" when (addr =  x"ad") else
x"0002" when (addr =  x"ae") else
x"0002" when (addr =  x"af") else
x"002D" when (addr =  x"b0") else
x"000A" when (addr =  x"b1") else
x"0002" when (addr =  x"b2") else
x"0002" when (addr =  x"b3") else
x"002D" when (addr =  x"b4") else
x"000A" when (addr =  x"b5") else
x"0002" when (addr =  x"b6") else
x"000A" when (addr =  x"b7") else
x"004C" when (addr =  x"b8") else
x"000A" when (addr =  x"b9") else
x"004C" when (addr =  x"ba") else
x"0002" when (addr =  x"bb") else
x"004D" when (addr =  x"bc") else
x"000A" when (addr =  x"bd") else
x"0002" when (addr =  x"be") else
x"0002" when (addr =  x"bf") else
x"004A" when (addr =  x"c0") else
x"000A" when (addr =  x"c1") else
x"0002" when (addr =  x"c2") else
x"0002" when (addr =  x"c3") else
x"005F" when (addr =  x"c4") else
x"000A" when (addr =  x"c5") else
x"0002" when (addr =  x"c6") else
x"0002" when (addr =  x"c7") else
x"0043" when (addr =  x"c8") else
x"000A" when (addr =  x"c9") else
x"0002" when (addr =  x"ca") else
x"0002" when (addr =  x"cb") else
x"0050" when (addr =  x"cc") else
x"000A" when (addr =  x"cd") else
x"0002" when (addr =  x"ce") else
x"0002" when (addr =  x"cf") else
x"0055" when (addr =  x"d0") else
x"000A" when (addr =  x"d1") else
x"0002" when (addr =  x"d2") else
x"0002" when (addr =  x"d3") else
x"0020" when (addr =  x"d4") else
x"000A" when (addr =  x"d5") else
x"0002" when (addr =  x"d6") else
x"0002" when (addr =  x"d7") else
x"004C" when (addr =  x"d8") else
x"000A" when (addr =  x"d9") else
x"0002" when (addr =  x"da") else
x"0002" when (addr =  x"db") else
x"006F" when (addr =  x"dc") else
x"000A" when (addr =  x"dd") else
x"0002" when (addr =  x"de") else
x"0002" when (addr =  x"df") else
x"0061" when (addr =  x"e0") else
x"000A" when (addr =  x"e1") else
x"0002" when (addr =  x"e2") else
x"0002" when (addr =  x"e3") else
x"0064" when (addr =  x"e4") else
x"000A" when (addr =  x"e5") else
x"0002" when (addr =  x"e6") else
x"0002" when (addr =  x"e7") else
x"0065" when (addr =  x"e8") else
x"000A" when (addr =  x"e9") else
x"0002" when (addr =  x"ea") else
x"0002" when (addr =  x"eb") else
x"0072" when (addr =  x"ec") else
x"000A" when (addr =  x"ed") else
x"0002" when (addr =  x"ee") else
x"0002" when (addr =  x"ef") else
x"0020" when (addr =  x"f0") else
x"000A" when (addr =  x"f1") else
x"0002" when (addr =  x"f2") else
x"0002" when (addr =  x"f3") else
x"0032" when (addr =  x"f4") else
x"000A" when (addr =  x"f5") else
x"0002" when (addr =  x"f6") else
x"0002" when (addr =  x"f7") else
x"002E" when (addr =  x"f8") else
x"000A" when (addr =  x"f9") else
x"0002" when (addr =  x"fa") else
x"0002" when (addr =  x"fb") else
x"0030" when (addr =  x"fc") else
x"000A" when (addr =  x"fd") else
x"0002" when (addr =  x"fe") else
x"0002" when (addr =  x"ff") else
x"000D" when (addr =  x"100") else
x"000A" when (addr =  x"101") else
x"0002" when (addr =  x"102") else
x"0002" when (addr =  x"103") else
x"000A" when (addr =  x"104") else
x"000A" when (addr =  x"105") else
x"0002" when (addr =  x"106") else
x"000A" when (addr =  x"107") else
x"004C" when (addr =  x"108") else
x"0002" when (addr =  x"109") else
x"002D" when (addr =  x"10a") else
x"000A" when (addr =  x"10b") else
x"0002" when (addr =  x"10c") else
x"0002" when (addr =  x"10d") else
x"002D" when (addr =  x"10e") else
x"000A" when (addr =  x"10f") else
x"0002" when (addr =  x"110") else
x"0002" when (addr =  x"111") else
x"002D" when (addr =  x"112") else
x"000A" when (addr =  x"113") else
x"0002" when (addr =  x"114") else
x"0002" when (addr =  x"115") else
x"002D" when (addr =  x"116") else
x"000A" when (addr =  x"117") else
x"0002" when (addr =  x"118") else
x"0002" when (addr =  x"119") else
x"002D" when (addr =  x"11a") else
x"000A" when (addr =  x"11b") else
x"0002" when (addr =  x"11c") else
x"0002" when (addr =  x"11d") else
x"002D" when (addr =  x"11e") else
x"000A" when (addr =  x"11f") else
x"0002" when (addr =  x"120") else
x"0002" when (addr =  x"121") else
x"002D" when (addr =  x"122") else
x"000A" when (addr =  x"123") else
x"0002" when (addr =  x"124") else
x"0002" when (addr =  x"125") else
x"002D" when (addr =  x"126") else
x"000A" when (addr =  x"127") else
x"0002" when (addr =  x"128") else
x"0002" when (addr =  x"129") else
x"002D" when (addr =  x"12a") else
x"000A" when (addr =  x"12b") else
x"0002" when (addr =  x"12c") else
x"0002" when (addr =  x"12d") else
x"002D" when (addr =  x"12e") else
x"000A" when (addr =  x"12f") else
x"0002" when (addr =  x"130") else
x"0002" when (addr =  x"131") else
x"002D" when (addr =  x"132") else
x"000A" when (addr =  x"133") else
x"0002" when (addr =  x"134") else
x"0002" when (addr =  x"135") else
x"002D" when (addr =  x"136") else
x"000A" when (addr =  x"137") else
x"0002" when (addr =  x"138") else
x"0002" when (addr =  x"139") else
x"002D" when (addr =  x"13a") else
x"000A" when (addr =  x"13b") else
x"0002" when (addr =  x"13c") else
x"0002" when (addr =  x"13d") else
x"002D" when (addr =  x"13e") else
x"000A" when (addr =  x"13f") else
x"0002" when (addr =  x"140") else
x"0002" when (addr =  x"141") else
x"002D" when (addr =  x"142") else
x"000A" when (addr =  x"143") else
x"0002" when (addr =  x"144") else
x"0002" when (addr =  x"145") else
x"002D" when (addr =  x"146") else
x"000A" when (addr =  x"147") else
x"0002" when (addr =  x"148") else
x"0002" when (addr =  x"149") else
x"002D" when (addr =  x"14a") else
x"000A" when (addr =  x"14b") else
x"0002" when (addr =  x"14c") else
x"000A" when (addr =  x"14d") else
x"004C" when (addr =  x"14e") else
x"000A" when (addr =  x"14f") else
x"004C" when (addr =  x"150") else
x"000A" when (addr =  x"151") else
x"0037" when (addr =  x"152") else
x"0002" when (addr =  x"153") else
x"0400" when (addr =  x"154") else
x"0008" when (addr =  x"155") else
x"000A" when (addr =  x"156") else
x"0037" when (addr =  x"157") else
x"0002" when (addr =  x"158") else
x"0401" when (addr =  x"159") else
x"0008" when (addr =  x"15a") else
x"0002" when (addr =  x"15b") else
x"0000" when (addr =  x"15c") else
x"0002" when (addr =  x"15d") else
x"0402" when (addr =  x"15e") else
x"0008" when (addr =  x"15f") else
x"0002" when (addr =  x"160") else
x"0402" when (addr =  x"161") else
x"0009" when (addr =  x"162") else
x"0002" when (addr =  x"163") else
x"0400" when (addr =  x"164") else
x"0009" when (addr =  x"165") else
x"0005" when (addr =  x"166") else
x"000C" when (addr =  x"167") else
x"017E" when (addr =  x"168") else
x"000A" when (addr =  x"169") else
x"0037" when (addr =  x"16a") else
x"0002" when (addr =  x"16b") else
x"0403" when (addr =  x"16c") else
--next line is no-op to fix a bug.
x"0001" when (addr =  x"16d") else
x"0002" when (addr =  x"16e") else
x"0402" when (addr =  x"16f") else
x"0009" when (addr =  x"170") else
x"0018" when (addr =  x"171") else
x"0008" when (addr =  x"172") else
x"0002" when (addr =  x"173") else
x"0402" when (addr =  x"174") else
x"0009" when (addr =  x"175") else
x"0002" when (addr =  x"176") else
x"0001" when (addr =  x"177") else
x"0018" when (addr =  x"178") else
x"0002" when (addr =  x"179") else
x"0402" when (addr =  x"17a") else
x"0008" when (addr =  x"17b") else
x"0004" when (addr =  x"17c") else
x"0160" when (addr =  x"17d") else
x"0002" when (addr =  x"17e") else
x"0401" when (addr =  x"17f") else
x"0009" when (addr =  x"180") else
x"000D" when (addr =  x"181") else
x"000B" when (addr =  x"182") else
x"0003"; -- Halt instruction 
      data <= output when cs = '0' else "ZZZZZZZZZZZZZZZZ";

end Behavioral;
